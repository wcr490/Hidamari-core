module peripheral_bus (
);
    
endmodule